module shiftreg